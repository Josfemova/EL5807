*Custom Compiler Version U-2023.03-SP2
*Wed Nov 27 23:46:34 2024

*.SCALE METER
*.LDD
.GLOBAL gnd! vdd!
********************************************************************************
* Library          : tarea2
* Cell             : nor2in
* View             : schematic
* View Search List : auCdl cmos_sch schematic
* View Stop List   : auCdl
********************************************************************************
.subckt nor2in A B Q
*.PININFO A:I B:I Q:O
MM3 Q B gnd! gnd! NE W=360n L=180n M='1*2' AD=9.72e-14 AS=1.728e-13 NRD=0.75
+ NRS=0.75 PD=9e-07 PS=1.68e-06
MM0 Q A gnd! gnd! NE W=360n L=180n M='1*2' AD=9.72e-14 AS=1.728e-13 NRD=0.75
+ NRS=0.75 PD=9e-07 PS=1.68e-06
MM2 Q B net9 vdd! PE W=720n L=180n M='1*4' AD=1.944e-13 AS=2.7e-13 NRD=0.375
+ NRS=0.375 PD=1.26e-06 PS=1.83e-06
MM1 net9 A vdd! vdd! PE W=720n L=180n M='1*4' AD=1.944e-13 AS=2.7e-13 NRD=0.375
+ NRS=0.375 PD=1.26e-06 PS=1.83e-06
.ends nor2in


