
.option post

.temp 70 
.param SUPPLY=1.8
.param H=4
.param N1=4
.param Ratio=2
.option scale=90n


.lib '/mnt/vol_NFS_rh003/Est_VLSI_II_2024/sfallas/EL5807/Tarea_1/Hspice/lpmos/xh018.lib' tm
.lib '/mnt/vol_NFS_rh003/Est_VLSI_II_2024/sfallas/EL5807/Tarea_1/Hspice/lpmos/param.lib' 3s
.lib '/mnt/vol_NFS_rh003/Est_VLSI_II_2024/sfallas/EL5807/Tarea_1/Hspice/lpmos/config.lib' default


.global vdd! gnd!


.subckt inv in out N=4 P=8
xm0 out in gnd! gnd! ne w='N' l=2
+ as='N*5' ad='N*5' ps='2*N+10' pd='2*N+10'
xm1 out in vdd! vdd! pe w='P' l=2
+ as='P*5' ad='P*5' ps='2*P+10' pd='2*P+10'
.ends inv



*----------------------------------------------------------------------
* Simulation netlist
*----------------------------------------------------------------------
Vdd vdd! gnd! 'SUPPLY'
Vin a gnd! PULSE 0 'SUPPLY' 0ps 100ps 100ps 900ps 2ns
X1 a b inv P='P1' * shape input waveform
X2 b c inv P='P1' M=4 * reshape input waveform
X3 c d inv P='P1' M=16 * device under test
X4 d e inv P='P1' M=64 * load
X5 e f inv P='P1' M=256 * load on load
*----------------------------------------------------------------------
* Optimization setup
*----------------------------------------------------------------------
.param P1=optrange(8,4,16) * search from 4 to 16, guess 8
.model optmod opt itropt=30 * maximum of 30 iterations
.measure bestratio param='P1/4' * compute best P/N ratio
*----------------------------------------------------------------------
* Stimulus
*----------------------------------------------------------------------
.tran 1ps 2ns SWEEP OPTIMIZE=optrange RESULTS=diff MODEL=optmod

.measure tpdr * rising propagation delay
+ TRIG v(c) VAL='SUPPLY/2' FALL=1 
+ TARG v(d) VAL='SUPPLY/2' RISE=1
.measure tpdf * falling propagation delay
+ TRIG v(c) VAL='SUPPLY/2' RISE=1
+ TARG v(d) VAL='SUPPLY/2' FALL=1 
.measure tpd param='(tpdr+tpdf)/2' goal=0 * average prop delay
.measure diff param='tpdr-tpdf' goal=0 * diff between delays

.option measform=1
.option numdgt=6

.end
