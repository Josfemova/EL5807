* SPICE	Wed Nov 27 02:39:16 2024	not1out
* icv_netlist Version RHEL64 U-2022.12-SP4.9133772 2023/08/28

* Hierarchy Level 0

* Top of hierarchy  cell=not1out
.subckt not1out gnd! vdd! Q A
X1 Q A gnd! gnd! ne  l=1.8e-07 w=3.6e-07 nrd=-1 nrs=-1 pd=1.88e-06 ps=1.04e-06
+	 ad=2.124e-13 as=1.242e-13
X2 gnd! A Q gnd! ne  l=1.8e-07 w=3.6e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.04e-06
+	 ad=1.242e-13 as=1.242e-13
X3 Q A gnd! gnd! ne  l=1.8e-07 w=3.6e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.04e-06
+	 ad=1.242e-13 as=1.242e-13
X4 gnd! A Q gnd! ne  l=1.8e-07 w=3.6e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.04e-06
+	 ad=1.242e-13 as=1.242e-13
X5 Q A gnd! gnd! ne  l=1.8e-07 w=3.6e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.04e-06
+	 ad=1.242e-13 as=1.242e-13
X6 gnd! A Q gnd! ne  l=1.8e-07 w=3.6e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.04e-06
+	 ad=1.242e-13 as=1.242e-13
X7 Q A gnd! gnd! ne  l=1.8e-07 w=3.6e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=3.62e-06
+	 ad=1.242e-13 as=5.448e-13
X8 gnd! vdd! p_dnw  area=3.05208e-11 pj=2.572e-05 perimeter=2.572e-05
X9 Q A vdd! vdd! pe  l=1.8e-07 w=7.2e-07 nrd=-1 nrs=-1 pd=2.4e-06 ps=1.26e-06
+	 ad=3.456e-13 as=1.944e-13
X10 vdd! A Q vdd! pe  l=1.8e-07 w=7.2e-07 nrd=-1 nrs=-1 pd=1.26e-06 ps=1.26e-06
+	 ad=1.944e-13 as=1.944e-13
X11 Q A vdd! vdd! pe  l=1.8e-07 w=7.2e-07 nrd=-1 nrs=-1 pd=1.26e-06 ps=1.26e-06
+	 ad=1.944e-13 as=1.944e-13
X12 vdd! A Q vdd! pe  l=1.8e-07 w=7.2e-07 nrd=-1 nrs=-1 pd=1.26e-06 ps=1.26e-06
+	 ad=1.944e-13 as=1.944e-13
X13 Q A vdd! vdd! pe  l=1.8e-07 w=7.2e-07 nrd=-1 nrs=-1 pd=1.26e-06 ps=1.26e-06
+	 ad=1.944e-13 as=1.944e-13
X14 vdd! A Q vdd! pe  l=1.8e-07 w=7.2e-07 nrd=-1 nrs=-1 pd=1.26e-06 ps=1.26e-06
+	 ad=1.944e-13 as=1.944e-13
X15 Q A vdd! vdd! pe  l=1.8e-07 w=7.2e-07 nrd=-1 nrs=-1 pd=1.26e-06 ps=5.04e-06
+	 ad=1.944e-13 as=7.108e-13
.ends not1out
